/***???????***/
module Pipeline_Control(Instruct,PC_sv,JT,Imm16,Shamt,Rd,Rt,Rs,PCSrc,RegDst,
  RegWr,ALUSrc1,ALUSrc2,ALUFun,Sign,MemWr,MemRd,MemToReg,EXTOp,LUOp,IRQ);
  
  input [31:0] Instruct;
  input PC_sv;
  output [25:0] JT;
  output [15:0] Imm16;
  output [4:0] Shamt,Rd,Rt,Rs;
  output [2:0] PCSrc;
  output [1:0] RegDst,MemToReg;
  output [5:0] ALUFun;
  output RegWr,ALUSrc1,ALUSrc2,Sign,MemWr,MemRd,EXTOp,LUOp;
  input IRQ;  //????
  
  wire  [5:0] Opcode, Funct;  //???????
  wire R,I,J,JR,nop;          //??????R?(JR??R???????)?J??I??????
  wire branch_con,branch_slt; //???????slt????
  wire normal;               //???????????????
  wire ILLOP,XADR;            //??????(ILLOP)????(XADR)

/*--------------------------------------------------------------------------*/
  
  assign Opcode=Instruct[31:26];//?????
  assign Funct=Instruct[5:0];   //??????????R?????
  
  assign JT=Instruct[25:0];     //target J?????
  assign Imm16=Instruct[15:0];  //??? I?????
  assign Shamt=Instruct[10:6];  //???R?????
  assign Rd=Instruct[15:11];    //R?????
  assign Rt=Instruct[20:16];    //R??I?????
  assign Rs=Instruct[25:21];    //R??I?????
 
  /*R?????add,addu,sub,subu,and,or,xor,nor,sll,srl,sra,jr,jalr?????R?1*/ 
  assign R= ~nop&(Opcode==6'b0)&
   			( (Instruct[10:3]==8'b00000100) |      //??add,addu,sub,subu,and,or,xor,nor ??
				(Instruct[10:0]==11'b00000101010) |  //??slt??
				((Instruct[25:21] == 5'd0)&(Instruct[5:2]==4'd0)&(Instruct[1:0]!=2'b01))| //??sll,srl,sra????
				({Instruct[20:11],Instruct[5:1]}==15'b000000000000100) |               //??jr??
				({Instruct[20:16],Instruct[5:0]}==11'b00000001001)                     //??jalr??
			);    
	
	/*I?????addi,addiu,andi,slti,sltiu,lui,lw,sw,beq,bne,blez,bgtz,bltz?????I?1*/
  assign I=
      ( ((Instruct[31:29]==3'b001)&((Instruct[28:26]==3'b100)|~Instruct[28]|(Instruct[28:21]==8'b11100000)))|  //????addi,addiu,andi,slti,sltiu,lui
			  ((Instruct[31:30]==2'b10)&(Instruct[28:26]==3'b011))|  //??lw,sw??
			  ((Instruct[31:29]==3'b000)&((Instruct[28:27]==2'b10)|  //??beq,bne??
			  ((Instruct[20:16]==5'b00000)&((Instruct[28:27]==2'b11)|(Instruct[28:26]==3'b001)))))//??blez,bgtz,bltz??
		  );
		  
	/*J???*/
	assign J=(Instruct[31:27]==5'b00001);  //??j,jal???????J?1
	/*R?????????*/	
	assign JR=R&(Instruct[5:1]==5'b00100); //??jr, jalr????
  /*??? nop (0x00000000,?sll $0,$0,0)*/
	assign nop=(Instruct==32'h0);  //????nop?1
	
  assign branch_con=I&(Instruct[31:29]==3'b000);  //????beq,bne,blez,bgtz,bltz????????branch_con=1
  assign branch_slt=(R&Instruct[3])|(I&~Instruct[31]
                  &(Instruct[28:27]==2'b01)); //????????slt,slti,sltiu??branch_slt=1
  assign normal=R|I|J|nop;   //R?I?J?nop????????????MIPS???????????????
  assign ILLOP=~PC_sv&IRQ;     //????0????????ILLOP=1
  assign XADR=~PC_sv&~normal;  //????0????????XADR=1
 
/*-----------------------------------------------------------------------------*/
 
/*???????*/
  //PCSrc
    /*???????????PCSc=001????????branch_con=1;
      PCSc=011?jr,jalr??,JR=1;PCSc=101????,XADR=1*/
    assign PCSrc[0]=(JR|branch_con|XADR)&~ILLOP;  
    /*???????????PCSrc=010????J=1?JR=1*/
    assign PCSrc[1]=(JR|J)&~ILLOP;
    /*PRSrc=100?101????????????*/
    assign PCSrc[2]=XADR|ILLOP;
    
  //RegDst:
    /*?????????RegDst=01????????Rt,??I???;
      RegDst=11????????Xp,?????????????????$26????*/
    assign RegDst[0]=I|~normal|XADR;//?
    /*?????????RegDst=10????????$ra??$31???;
      RegDst=11????????Xp,?????????????????$26????*/
    assign RegDst[1]=MemToReg[1]|~normal;//?
   
  //RegWr
  /*??????????R??Jr??(??31????)?jal???I?????addi,addiu,andi,
    slti,sltiu,lui????????????26????????????RegWr???1*/
    assign RegWr=(R&~(JR&~Funct[0]))|(I&~branch_con&~MemWr)|(J&Opcode[0])|XADR;
    
  //ALUSrc1
  /*ALUSrc1=1?,??shamt[4:0],????????,sll,srl,sra?Funct[5:0]??
    ???000000?000010?000100?add?addu?and?sub?subu?or?nor?xor?Funct[5]??1,
    jr?jalr?Funct[5]??0??Funct[3]??1*/
    assign ALUSrc1=R&~Funct[5]&~Funct[3];  //sll,srl,sra
  
  //ALUSrc2
  /*ALUSrc2=1??????????????????I?????????????*/
    assign ALUSrc2=I&~branch_con; 
    
  //ALUFun
    /*ALUFun=[5:4]=00?,???????;01????????;10???????;11??????*/
    assign ALUFun[5]=(R&~Funct[5])|branch_con|branch_slt; //??????j??               
    assign ALUFun[4]=(R&Funct[2])|branch_con|branch_slt|(Opcode[3:1]==3'b110); //???????
    /*(R&(Funct[2:1]==2'b10))??and?or;(branch_con&Opcode[1])??blez,bgtz??;
      (Opcode[3:1]==3'b110)??andi??*/
    assign ALUFun[3]=(R&(Funct[2:1]==2'b10))|(branch_con&Opcode[1])|(Opcode[3:1]==3'b110); //??and,or,blez,bgtz,andi??
    assign ALUFun[2]=(R&Funct[2]&(Funct[1]^Funct[0]))|((branch_con|branch_slt)&(Opcode[2:1]!=2'b10));//??or,xor,bgtz,blez,bltz,slt,slti,sltiu??
    assign ALUFun[1]=(R&Funct[2]&(Funct[1]^Funct[0]))|(R&Funct[0]&~Funct[5])|
                    (((Opcode[2:0]==3'b100)|(Opcode[2:0]==3'b111))&branch_con); //??or,xor,sra,jalr,beq,bgtz??
    assign ALUFun[0]=(R&Funct[1]&(~Funct[2]|Funct[0]))|branch_con|branch_slt; //??sub,subi,nor,srl,sra,slt??
  
  //Sign
    /*Sign??ALU??????????????????Sign=1????????
      ??R????and,sub?I????addi,slt*/                 
    assign Sign=(R&(Funct[5:2]==4'b1000)&~Funct[0])|(I&(Opcode[5:2]==4'b0010)&~Opcode[0]);
    
  //MemRd
    /*?????????lw??*/
    assign MemRd=Opcode[5]&~Opcode[3]; //Opcode==6'b100011
    
  //MemWr
    /*?????????sw??*/
    assign MemWr=Opcode[5]&Opcode[3];  //Opcode==6'b101011
  
  //MemToReg
    /*??????????????MemToReg=00????ALU?????;
      MemToReg=01???????????????lw??;MemToReg=10????PC+4*/
    assign MemToReg[0]=MemRd;  
    assign MemToReg[1]=(J&Opcode[0])|(JR&Funct[0])|XADR; /*????jal?jalr?????*/
    
  //EXTOp
    /*EXTOp???????16?????32????????????????
      EXTOp=1???????*/
    assign EXTOp=Sign;
    
  //LUOp
    /*????lui??16??????32????16??*/
    assign LUOp=(Opcode[3:1]==3'b111); //lui
endmodule

