module seqdetector_Reg(clk_in,system_clk,reset,x,z,leds);
  input clk_in,system_clk,reset,x;//?????system_clk?????????????clk_in??????reset??????x???
  output reg z;//????
  output reg [6:1] leds;//?????????6?LED??
  wire clk_o;//????????????
  
  debounce d(system_clk,clk_in,clk_o);//????
  
  always @(posedge clk_o or posedge reset)
    begin
      if(reset) 
        leds<=0;//???????????
      else 
      begin
        leds=(leds<<1);//?????
        leds[1]=x;//??????????
      end
    end
  
  always @(leds)//???????????????
    begin
      if(leds==6'b101011) z<=1;//??????????????1
      else z<=0;
    end
endmodule
