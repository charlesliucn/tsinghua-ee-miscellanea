/*?100MHz??????1Hz??????*/
module gen_clk(sysclk,clk_ctrl,clk_scan); 
  input sysclk; 
  output reg clk_ctrl,clk_scan; 
  reg [31:0]count1;//100MHz?????100000000??????1Hz?????1???
  reg [31:0]count2;//100MHz?????100000??????1kHz?????1???
  initial//???
  begin 
    clk_ctrl<=0;
    clk_scan<=0; 
    count1<=0;
    count2<=0;
  end 
  always@(posedge sysclk)//??????????? 
  begin 
  if(count1==32'd49999999) 
    begin 
      clk_ctrl<=~clk_ctrl; 
      count1<=0; 
    end 
  else 
    count1<=count1+32'd1;
  end
  always@(posedge sysclk)//??????????? 
  begin 
  if(count2==32'd49999) 
    begin 
      clk_scan<=~clk_scan; 
      count2<=0; 
    end 
  else 
    count2<=count2+32'd1;
  end
endmodule
