module synaddcounter(leds,ano,btnd,reset,clk);
output [6:0]leds;//??led?7????
output [3:0]ano;//??????LED????
input btnd,reset,clk;//btnd????????
reg [3:0]Q;//?????
wire BTND;//BTND?????????????

assign ano=4'b0000;//4?LED??
debounce d(clk,btnd,BTND);//????
always @(posedge BTND or posedge reset)//???????????????
  begin
  if(reset) //???0
    begin 
      Q[1]<=0;
      Q[2]<=0;
      Q[3]<=0;
      Q[0]<=0; 
  end
  else //????
    begin
      Q[0]<=~Q[0];
      if(Q[0]) 
      begin
        Q[1]<=~Q[1];
        if(Q[1]) 
        begin
          Q[2]<=~Q[2];
          if(Q[2]) 
          begin
            Q[3]<=~Q[3];
          end
        end
      end
    end
  end
BCD7 bcd7(Q,leds);
endmodule

