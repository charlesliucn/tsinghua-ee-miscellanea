module spanmode(modecontrol,sigin,sigout);
  input sigin,modecontrol;//???????????
  output sigout; //????
  reg sigout_temp;
  reg [3:0]count; //?????????
  assign sigout=sigout_temp;
  initial
    begin
      sigout_temp<=0; //???
      count<=0; 
    end

  always @(posedge sigin)//???????????
    begin 
      if(~modecontrol)//modecontrol????????????
        sigout_temp=~sigout_temp;
      else//modecontrol??????????????????????
        begin 
          if(count==4) 
            begin 
              sigout_temp<=~sigout_temp; 
              count<=0; 
            end
          else 
            count<=count+1; 
        end 
    end
endmodule
