/*指令存储器单元*/
module CPU_ROM(addr,data);
  input [6:0] addr;
  output reg[31:0] data;
  
  always@(*) 
  begin
		case(addr[6:0])
		7'd0:data<=32'b00001000000000000000000001001010;
        7'd1:data<=32'b00001000000000000000000001010000;
        7'd2:data<=32'b00000011010000000000000000001000;
        7'd3:data<=32'b00100100000001000000000011000000;
        7'd4:data<=32'b10101100000001000000000000000000;
        7'd5:data<=32'b00100100000001000000000011111001;
        7'd6:data<=32'b10101100000001000000000000000100;
        7'd7:data<=32'b00100100000001000000000010100100;
        7'd8:data<=32'b10101100000001000000000000001000;
        7'd9:data<=32'b00100100000001000000000010110000;
        7'd10:data<=32'b10101100000001000000000000001100;
        7'd11:data<=32'b00100100000001000000000010011001;
        7'd12:data<=32'b10101100000001000000000000010000;
        7'd13:data<=32'b00100100000001000000000010010010;
        7'd14:data<=32'b10101100000001000000000000010100;
        7'd15:data<=32'b00100100000001000000000010000010;
        7'd16:data<=32'b10101100000001000000000000011000;
        7'd17:data<=32'b00100100000001000000000011111000;
        7'd18:data<=32'b10101100000001000000000000011100;
        7'd19:data<=32'b00100100000001000000000010000000;
        7'd20:data<=32'b10101100000001000000000000100000;
        7'd21:data<=32'b00100100000001000000000010010000;
        7'd22:data<=32'b10101100000001000000000000100100;
        7'd23:data<=32'b00100100000001000000000010001000;
        7'd24:data<=32'b10101100000001000000000000101000;
        7'd25:data<=32'b00100100000001000000000010000011;
        7'd26:data<=32'b10101100000001000000000000101100;
        7'd27:data<=32'b00100100000001000000000011000110;
        7'd28:data<=32'b10101100000001000000000000110000;
        7'd29:data<=32'b00100100000001000000000010100001;
        7'd30:data<=32'b10101100000001000000000000110100;
        7'd31:data<=32'b00100100000001000000000010000110;
        7'd32:data<=32'b10101100000001000000000000111000;
        7'd33:data<=32'b00100100000001000000000010001110;
        7'd34:data<=32'b10101100000001000000000000111100;
        7'd35:data<=32'b00100100000000100000000000000001;
        7'd36:data<=32'b10001110000100010000000000011100;
        7'd37:data<=32'b00000010001000000010100000100000;
        7'd38:data<=32'b10001110000100100000000000011100;
        7'd39:data<=32'b00000010010000000011000000100000;
        7'd40:data<=32'b00010000000001010000000000001000;
        7'd41:data<=32'b00010000000001100000000000001001;
        7'd42:data<=32'b00010000110001010000000000001000;
        7'd43:data<=32'b00000000101001100010000000101010;
        7'd44:data<=32'b00010100000001000000000000000010;
        7'd45:data<=32'b00000000101001100010100000100010;
        7'd46:data<=32'b00001000000000000000000000101010;
        7'd47:data<=32'b00000000110001010011000000100010;
        7'd48:data<=32'b00001000000000000000000000101010;
        7'd49:data<=32'b00000000110000000001100000100000;
        7'd50:data<=32'b00001000000000000000000000110100;
        7'd51:data<=32'b00000000101000000001100000100000;
        7'd52:data<=32'b00000000000000100100000001000010;
        7'd53:data<=32'b00010000000010000000000000001000;
        7'd54:data<=32'b00000000000000100100000010000010;
        7'd55:data<=32'b00010000000010000000000000001001;
        7'd56:data<=32'b00000000000000100100000011000010;
        7'd57:data<=32'b00010000000010000000000000001010;
        7'd58:data<=32'b00100100000000100000000000000001;
        7'd59:data<=32'b00110010001100110000000000001111;
        7'd60:data<=32'b00000000000100111001100010000000;
        7'd61:data<=32'b00001000000000000000000001001000;
        7'd62:data<=32'b00000000000100011001100100000010;
        7'd63:data<=32'b00000000000100111001100010000000;
        7'd64:data<=32'b00001000000000000000000001000111;
        7'd65:data<=32'b00110010010100110000000000001111;
        7'd66:data<=32'b00000000000100111001100010000000;
        7'd67:data<=32'b00001000000000000000000001000111;
        7'd68:data<=32'b00000000000100101001100100000010;
        7'd69:data<=32'b00000000000100111001100010000000;
        7'd70:data<=32'b00001000000000000000000001000111;
        7'd71:data<=32'b00000000000000100001000001000000;
        7'd72:data<=32'b00001000000000000000000001001000;
        7'd73:data<=32'b00001000000000000000000000100100;
        7'd74:data<=32'b00100100000101000000000000000011;
        7'd75:data<=32'b00111100000100000100000000000000;
        7'd76:data<=32'b10101110000101000000000000001000;
        7'd77:data<=32'b00100100000101110000000000000011;
        7'd78:data<=32'b00000000000101111011100010000000;
        7'd79:data<=32'b00000010111000000000000000001000;
        7'd80:data<=32'b10101110000101000000000000001000;
        7'd81:data<=32'b10001110011101010000000000000000;
        7'd82:data<=32'b00000000000000101011001000000000;
        7'd83:data<=32'b00000010101101101011000000100000;
        7'd84:data<=32'b10101110000101100000000000010100;
        7'd85:data<=32'b10101110000000110000000000001100;
        7'd86:data<=32'b10101110000000110000000000011000;
        7'd87:data<=32'b00000011111000000000000000001000;
		 default:	data<=32'b0;
		endcase
 end
endmodule